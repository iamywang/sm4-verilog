module sbox (input [7:0] data_in,
             output reg [7:0] res_out);

always@(*)
    case(data_in)
        8'h00 : res_out <= 8'hd6;
        8'h01 : res_out <= 8'h90;
        8'h02 : res_out <= 8'he9;
        8'h03 : res_out <= 8'hfe;
        8'h04 : res_out <= 8'hcc;
        8'h05 : res_out <= 8'he1;
        8'h06 : res_out <= 8'h3d;
        8'h07 : res_out <= 8'hb7;
        8'h08 : res_out <= 8'h16;
        8'h09 : res_out <= 8'hb6;
        8'h0a : res_out <= 8'h14;
        8'h0b : res_out <= 8'hc2;
        8'h0c : res_out <= 8'h28;
        8'h0d : res_out <= 8'hfb;
        8'h0e : res_out <= 8'h2c;
        8'h0f : res_out <= 8'h05;
        8'h10 : res_out <= 8'h2b;
        8'h11 : res_out <= 8'h67;
        8'h12 : res_out <= 8'h9a;
        8'h13 : res_out <= 8'h76;
        8'h14 : res_out <= 8'h2a;
        8'h15 : res_out <= 8'hbe;
        8'h16 : res_out <= 8'h04;
        8'h17 : res_out <= 8'hc3;
        8'h18 : res_out <= 8'haa;
        8'h19 : res_out <= 8'h44;
        8'h1a : res_out <= 8'h13;
        8'h1b : res_out <= 8'h26;
        8'h1c : res_out <= 8'h49;
        8'h1d : res_out <= 8'h86;
        8'h1e : res_out <= 8'h06;
        8'h1f : res_out <= 8'h99;
        8'h20 : res_out <= 8'h9c;
        8'h21 : res_out <= 8'h42;
        8'h22 : res_out <= 8'h50;
        8'h23 : res_out <= 8'hf4;
        8'h24 : res_out <= 8'h91;
        8'h25 : res_out <= 8'hef;
        8'h26 : res_out <= 8'h98;
        8'h27 : res_out <= 8'h7a;
        8'h28 : res_out <= 8'h33;
        8'h29 : res_out <= 8'h54;
        8'h2a : res_out <= 8'h0b;
        8'h2b : res_out <= 8'h43;
        8'h2c : res_out <= 8'hed;
        8'h2d : res_out <= 8'hcf;
        8'h2e : res_out <= 8'hac;
        8'h2f : res_out <= 8'h62;
        8'h30 : res_out <= 8'he4;
        8'h31 : res_out <= 8'hb3;
        8'h32 : res_out <= 8'h1c;
        8'h33 : res_out <= 8'ha9;
        8'h34 : res_out <= 8'hc9;
        8'h35 : res_out <= 8'h08;
        8'h36 : res_out <= 8'he8;
        8'h37 : res_out <= 8'h95;
        8'h38 : res_out <= 8'h80;
        8'h39 : res_out <= 8'hdf;
        8'h3a : res_out <= 8'h94;
        8'h3b : res_out <= 8'hfa;
        8'h3c : res_out <= 8'h75;
        8'h3d : res_out <= 8'h8f;
        8'h3e : res_out <= 8'h3f;
        8'h3f : res_out <= 8'ha6;
        8'h40 : res_out <= 8'h47;
        8'h41 : res_out <= 8'h07;
        8'h42 : res_out <= 8'ha7;
        8'h43 : res_out <= 8'hfc;
        8'h44 : res_out <= 8'hf3;
        8'h45 : res_out <= 8'h73;
        8'h46 : res_out <= 8'h17;
        8'h47 : res_out <= 8'hba;
        8'h48 : res_out <= 8'h83;
        8'h49 : res_out <= 8'h59;
        8'h4a : res_out <= 8'h3c;
        8'h4b : res_out <= 8'h19;
        8'h4c : res_out <= 8'he6;
        8'h4d : res_out <= 8'h85;
        8'h4e : res_out <= 8'h4f;
        8'h4f : res_out <= 8'ha8;
        8'h50 : res_out <= 8'h68;
        8'h51 : res_out <= 8'h6b;
        8'h52 : res_out <= 8'h81;
        8'h53 : res_out <= 8'hb2;
        8'h54 : res_out <= 8'h71;
        8'h55 : res_out <= 8'h64;
        8'h56 : res_out <= 8'hda;
        8'h57 : res_out <= 8'h8b;
        8'h58 : res_out <= 8'hf8;
        8'h59 : res_out <= 8'heb;
        8'h5a : res_out <= 8'h0f;
        8'h5b : res_out <= 8'h4b;
        8'h5c : res_out <= 8'h70;
        8'h5d : res_out <= 8'h56;
        8'h5e : res_out <= 8'h9d;
        8'h5f : res_out <= 8'h35;
        8'h60 : res_out <= 8'h1e;
        8'h61 : res_out <= 8'h24;
        8'h62 : res_out <= 8'h0e;
        8'h63 : res_out <= 8'h5e;
        8'h64 : res_out <= 8'h63;
        8'h65 : res_out <= 8'h58;
        8'h66 : res_out <= 8'hd1;
        8'h67 : res_out <= 8'ha2;
        8'h68 : res_out <= 8'h25;
        8'h69 : res_out <= 8'h22;
        8'h6a : res_out <= 8'h7c;
        8'h6b : res_out <= 8'h3b;
        8'h6c : res_out <= 8'h01;
        8'h6d : res_out <= 8'h21;
        8'h6e : res_out <= 8'h78;
        8'h6f : res_out <= 8'h87;
        8'h70 : res_out <= 8'hd4;
        8'h71 : res_out <= 8'h00;
        8'h72 : res_out <= 8'h46;
        8'h73 : res_out <= 8'h57;
        8'h74 : res_out <= 8'h9f;
        8'h75 : res_out <= 8'hd3;
        8'h76 : res_out <= 8'h27;
        8'h77 : res_out <= 8'h52;
        8'h78 : res_out <= 8'h4c;
        8'h79 : res_out <= 8'h36;
        8'h7a : res_out <= 8'h02;
        8'h7b : res_out <= 8'he7;
        8'h7c : res_out <= 8'ha0;
        8'h7d : res_out <= 8'hc4;
        8'h7e : res_out <= 8'hc8;
        8'h7f : res_out <= 8'h9e;
        8'h80 : res_out <= 8'hea;
        8'h81 : res_out <= 8'hbf;
        8'h82 : res_out <= 8'h8a;
        8'h83 : res_out <= 8'hd2;
        8'h84 : res_out <= 8'h40;
        8'h85 : res_out <= 8'hc7;
        8'h86 : res_out <= 8'h38;
        8'h87 : res_out <= 8'hb5;
        8'h88 : res_out <= 8'ha3;
        8'h89 : res_out <= 8'hf7;
        8'h8a : res_out <= 8'hf2;
        8'h8b : res_out <= 8'hce;
        8'h8c : res_out <= 8'hf9;
        8'h8d : res_out <= 8'h61;
        8'h8e : res_out <= 8'h15;
        8'h8f : res_out <= 8'ha1;
        8'h90 : res_out <= 8'he0;
        8'h91 : res_out <= 8'hae;
        8'h92 : res_out <= 8'h5d;
        8'h93 : res_out <= 8'ha4;
        8'h94 : res_out <= 8'h9b;
        8'h95 : res_out <= 8'h34;
        8'h96 : res_out <= 8'h1a;
        8'h97 : res_out <= 8'h55;
        8'h98 : res_out <= 8'had;
        8'h99 : res_out <= 8'h93;
        8'h9a : res_out <= 8'h32;
        8'h9b : res_out <= 8'h30;
        8'h9c : res_out <= 8'hf5;
        8'h9d : res_out <= 8'h8c;
        8'h9e : res_out <= 8'hb1;
        8'h9f : res_out <= 8'he3;
        8'ha0 : res_out <= 8'h1d;
        8'ha1 : res_out <= 8'hf6;
        8'ha2 : res_out <= 8'he2;
        8'ha3 : res_out <= 8'h2e;
        8'ha4 : res_out <= 8'h82;
        8'ha5 : res_out <= 8'h66;
        8'ha6 : res_out <= 8'hca;
        8'ha7 : res_out <= 8'h60;
        8'ha8 : res_out <= 8'hc0;
        8'ha9 : res_out <= 8'h29;
        8'haa : res_out <= 8'h23;
        8'hab : res_out <= 8'hab;
        8'hac : res_out <= 8'h0d;
        8'had : res_out <= 8'h53;
        8'hae : res_out <= 8'h4e;
        8'haf : res_out <= 8'h6f;
        8'hb0 : res_out <= 8'hd5;
        8'hb1 : res_out <= 8'hdb;
        8'hb2 : res_out <= 8'h37;
        8'hb3 : res_out <= 8'h45;
        8'hb4 : res_out <= 8'hde;
        8'hb5 : res_out <= 8'hfd;
        8'hb6 : res_out <= 8'h8e;
        8'hb7 : res_out <= 8'h2f;
        8'hb8 : res_out <= 8'h03;
        8'hb9 : res_out <= 8'hff;
        8'hba : res_out <= 8'h6a;
        8'hbb : res_out <= 8'h72;
        8'hbc : res_out <= 8'h6d;
        8'hbd : res_out <= 8'h6c;
        8'hbe : res_out <= 8'h5b;
        8'hbf : res_out <= 8'h51;
        8'hc0 : res_out <= 8'h8d;
        8'hc1 : res_out <= 8'h1b;
        8'hc2 : res_out <= 8'haf;
        8'hc3 : res_out <= 8'h92;
        8'hc4 : res_out <= 8'hbb;
        8'hc5 : res_out <= 8'hdd;
        8'hc6 : res_out <= 8'hbc;
        8'hc7 : res_out <= 8'h7f;
        8'hc8 : res_out <= 8'h11;
        8'hc9 : res_out <= 8'hd9;
        8'hca : res_out <= 8'h5c;
        8'hcb : res_out <= 8'h41;
        8'hcc : res_out <= 8'h1f;
        8'hcd : res_out <= 8'h10;
        8'hce : res_out <= 8'h5a;
        8'hcf : res_out <= 8'hd8;
        8'hd0 : res_out <= 8'h0a;
        8'hd1 : res_out <= 8'hc1;
        8'hd2 : res_out <= 8'h31;
        8'hd3 : res_out <= 8'h88;
        8'hd4 : res_out <= 8'ha5;
        8'hd5 : res_out <= 8'hcd;
        8'hd6 : res_out <= 8'h7b;
        8'hd7 : res_out <= 8'hbd;
        8'hd8 : res_out <= 8'h2d;
        8'hd9 : res_out <= 8'h74;
        8'hda : res_out <= 8'hd0;
        8'hdb : res_out <= 8'h12;
        8'hdc : res_out <= 8'hb8;
        8'hdd : res_out <= 8'he5;
        8'hde : res_out <= 8'hb4;
        8'hdf : res_out <= 8'hb0;
        8'he0 : res_out <= 8'h89;
        8'he1 : res_out <= 8'h69;
        8'he2 : res_out <= 8'h97;
        8'he3 : res_out <= 8'h4a;
        8'he4 : res_out <= 8'h0c;
        8'he5 : res_out <= 8'h96;
        8'he6 : res_out <= 8'h77;
        8'he7 : res_out <= 8'h7e;
        8'he8 : res_out <= 8'h65;
        8'he9 : res_out <= 8'hb9;
        8'hea : res_out <= 8'hf1;
        8'heb : res_out <= 8'h09;
        8'hec : res_out <= 8'hc5;
        8'hed : res_out <= 8'h6e;
        8'hee : res_out <= 8'hc6;
        8'hef : res_out <= 8'h84;
        8'hf0 : res_out <= 8'h18;
        8'hf1 : res_out <= 8'hf0;
        8'hf2 : res_out <= 8'h7d;
        8'hf3 : res_out <= 8'hec;
        8'hf4 : res_out <= 8'h3a;
        8'hf5 : res_out <= 8'hdc;
        8'hf6 : res_out <= 8'h4d;
        8'hf7 : res_out <= 8'h20;
        8'hf8 : res_out <= 8'h79;
        8'hf9 : res_out <= 8'hee;
        8'hfa : res_out <= 8'h5f;
        8'hfb : res_out <= 8'h3e;
        8'hfc : res_out <= 8'hd7;
        8'hfd : res_out <= 8'hcb;
        8'hfe : res_out <= 8'h39;
        8'hff : res_out <= 8'h48;
    endcase

endmodule
